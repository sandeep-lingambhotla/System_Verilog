module test(a,b);
  
  input a;
  output b;
  
  assign #5 b = a;
  
endmodule
  
  
